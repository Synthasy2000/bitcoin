----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    01:53:54 06/02/2011
-- Design Name:
-- Module Name:    sha256_ch - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sha256_ch is
  Port ( x : in  STD_LOGIC_VECTOR (31 downto 0);
         y : in  STD_LOGIC_VECTOR (31 downto 0);
         z : in  STD_LOGIC_VECTOR (31 downto 0);
         q : out  STD_LOGIC_VECTOR (31 downto 0));
end sha256_ch;

architecture Behavioral of sha256_ch is

begin

  --listed in spec as: '(x and y) xor ((not x) and z)'
  --is 'z xor (x and (y xor z))' easier to implement in FPGA logic?
  q <= (x and y) xor ((not x) and z);

end Behavioral;

