----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    01:53:21 06/02/2011
-- Design Name:
-- Module Name:    sha256_e1 - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sha256_e1 is
  Port ( d : in  STD_LOGIC_VECTOR (31 downto 0);
         q : out  STD_LOGIC_VECTOR (31 downto 0));
end sha256_e1;

architecture Behavioral of sha256_e1 is

begin

  q <= (d(5 downto 0) & d(31 downto 6)) xor (d(10 downto 0) & d(31 downto 11)) xor (d(24 downto 0) & d(31 downto 25));

end Behavioral;

